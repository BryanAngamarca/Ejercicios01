----------------------------------------------------------------------------------
-- Create Date:    18:22:12 07/06/2022 
-- Module Name:    Rep_15 - Behavioral 
-- Bryan Angamarca
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Rep_15 is
    Port ( clk, reset : in  STD_LOGIC;
           q : inout  integer range 0 to 15);
end Replica_15_cont;

architecture Behavioral of Rep_15 is

begin
	process(clk, reset)
	begin
		if(clk' event and clk='1') then
			if(reset='1' or q=9) then
				q <= 0;
			else
				q <= q+1;
			end if;
		end if;
	end process;
end Behavioral;